LIBRARY IEEE;
USE STD.STANDARD.ALL;
ENTITY SUPER_CONTADOR IS
PORT( W,X,Y,Z: IN BIT;
		S: OUT BIT_VECTOR(3 DOWNTO 0));
		END SUPER_CONTADOR;
		
		
ARCHITECTURE CONTADOR OF SUPER_CONTADOR IS
SIGNAL ENTRADAS : BIT_VECTOR (3 DOWNTO 0);

BEGIN
ENTRADAS <= (W & X & Y & Z);

WITH ENTRADAS SELECT
	S <=  "0000" WHEN "0000",
	-- FULL 
			"0100" WHEN "1111",
			-- 3 
			"0011" WHEN "1110",
			"0011" WHEN "1101",
			"0011" WHEN "1011",
			"0011" WHEN "0111",
			-- 1 
			"0001" WHEN "0001",
			"0001" WHEN "0010",
			"0001" WHEN "0100",
			"0001" WHEN "1000",
			-- 2 
			"0010" WHEN OTHERS;
	
END CONTADOR;
			
			